`timescale 1ns / 1ps

module pol_mul_tb(

);

    reg [15:0] input_poly1;
	reg [15:0] input_poly2;
	
    reg start;
    reg clk, rst;
    wire [5:0] data_loop;
    
    wire [15:0] NTT_0, NTT_1, NTT_2, NTT_3, NTT_4, NTT_5, NTT_6, NTT_7, 
           NTT_8, NTT_9, NTT_10, NTT_11, NTT_12, NTT_13, NTT_14, NTT_15;
    
        
    wire [15:0] INTT_0, INTT_1, INTT_2, INTT_3, INTT_4, INTT_5, INTT_6, INTT_7, 
           INTT_8, INTT_9, INTT_10, INTT_11, INTT_12, INTT_13, INTT_14, INTT_15;
           
    Poly_mul dut(

            input_poly1, input_poly2, start, clk, rst, data_loop,
    
           NTT_0, NTT_1, NTT_2, NTT_3, NTT_4, NTT_5, NTT_6, NTT_7, 
           NTT_8, NTT_9, NTT_10, NTT_11, NTT_12, NTT_13, NTT_14, NTT_15,
      
           INTT_0, INTT_1, INTT_2, INTT_3, INTT_4, INTT_5, INTT_6, INTT_7, 
           INTT_8, INTT_9, INTT_10, INTT_11, INTT_12, INTT_13, INTT_14, INTT_15
    );
    
    initial
    begin
      clk = 1'b0; rst = 1'b0;
      forever #5 clk = ~clk;
    end
    
    initial
    begin
	#0 start = 1'b0; input_poly1 = 16'd257; input_poly2 = 16'd1;
	#10 start = 1'b1; input_poly1 = 16'd1; input_poly2 = 16'd257;
	#10 start = 1'b1; input_poly1 = 16'd2; input_poly2 = 16'd258;
	#10 start = 1'b1; input_poly1 = 16'd3; input_poly2 = 16'd259;
	#10 start = 1'b1; input_poly1 = 16'd4; input_poly2 = 16'd260;
	#10 start = 1'b1; input_poly1 = 16'd5; input_poly2 = 16'd261;
	#10 start = 1'b1; input_poly1 = 16'd6; input_poly2 = 16'd262;
	#10 start = 1'b1; input_poly1 = 16'd7; input_poly2 = 16'd263;
	#10 start = 1'b1; input_poly1 = 16'd8; input_poly2 = 16'd264;
	#10 start = 1'b1; input_poly1 = 16'd9; input_poly2 = 16'd265;
	#10 start = 1'b1; input_poly1 = 16'd10; input_poly2 = 16'd266;
	#10 start = 1'b1; input_poly1 = 16'd11; input_poly2 = 16'd267;
	#10 start = 1'b1; input_poly1 = 16'd12; input_poly2 = 16'd268;
	#10 start = 1'b1; input_poly1 = 16'd13; input_poly2 = 16'd269;
	#10 start = 1'b1; input_poly1 = 16'd14; input_poly2 = 16'd270;
	#10 start = 1'b1; input_poly1 = 16'd15; input_poly2 = 16'd271;
	#10 start = 1'b1; input_poly1 = 16'd16; input_poly2 = 16'd272;
	#10 start = 1'b1; input_poly1 = 16'd17; input_poly2 = 16'd273;
	#10 start = 1'b1; input_poly1 = 16'd18; input_poly2 = 16'd274;
	#10 start = 1'b1; input_poly1 = 16'd19; input_poly2 = 16'd275;
	#10 start = 1'b1; input_poly1 = 16'd20; input_poly2 = 16'd276;
	#10 start = 1'b1; input_poly1 = 16'd21; input_poly2 = 16'd277;
	#10 start = 1'b1; input_poly1 = 16'd22; input_poly2 = 16'd278;
	#10 start = 1'b1; input_poly1 = 16'd23; input_poly2 = 16'd279;
	#10 start = 1'b1; input_poly1 = 16'd24; input_poly2 = 16'd280;
	#10 start = 1'b1; input_poly1 = 16'd25; input_poly2 = 16'd281;
	#10 start = 1'b1; input_poly1 = 16'd26; input_poly2 = 16'd282;
	#10 start = 1'b1; input_poly1 = 16'd27; input_poly2 = 16'd283;
	#10 start = 1'b1; input_poly1 = 16'd28; input_poly2 = 16'd284;
	#10 start = 1'b1; input_poly1 = 16'd29; input_poly2 = 16'd285;
	#10 start = 1'b1; input_poly1 = 16'd30; input_poly2 = 16'd286;
	#10 start = 1'b1; input_poly1 = 16'd31; input_poly2 = 16'd287;
	#10 start = 1'b1; input_poly1 = 16'd32; input_poly2 = 16'd288;
	#10 start = 1'b1; input_poly1 = 16'd33; input_poly2 = 16'd289;
	#10 start = 1'b1; input_poly1 = 16'd34; input_poly2 = 16'd290;
	#10 start = 1'b1; input_poly1 = 16'd35; input_poly2 = 16'd291;
	#10 start = 1'b1; input_poly1 = 16'd36; input_poly2 = 16'd292;
	#10 start = 1'b1; input_poly1 = 16'd37; input_poly2 = 16'd293;
	#10 start = 1'b1; input_poly1 = 16'd38; input_poly2 = 16'd294;
	#10 start = 1'b1; input_poly1 = 16'd39; input_poly2 = 16'd295;
	#10 start = 1'b1; input_poly1 = 16'd40; input_poly2 = 16'd296;
	#10 start = 1'b1; input_poly1 = 16'd41; input_poly2 = 16'd297;
	#10 start = 1'b1; input_poly1 = 16'd42; input_poly2 = 16'd298;
	#10 start = 1'b1; input_poly1 = 16'd43; input_poly2 = 16'd299;
	#10 start = 1'b1; input_poly1 = 16'd44; input_poly2 = 16'd300;
	#10 start = 1'b1; input_poly1 = 16'd45; input_poly2 = 16'd301;
	#10 start = 1'b1; input_poly1 = 16'd46; input_poly2 = 16'd302;
	#10 start = 1'b1; input_poly1 = 16'd47; input_poly2 = 16'd303;
	#10 start = 1'b1; input_poly1 = 16'd48; input_poly2 = 16'd304;
	#10 start = 1'b1; input_poly1 = 16'd49; input_poly2 = 16'd305;
	#10 start = 1'b1; input_poly1 = 16'd50; input_poly2 = 16'd306;
	#10 start = 1'b1; input_poly1 = 16'd51; input_poly2 = 16'd307;
	#10 start = 1'b1; input_poly1 = 16'd52; input_poly2 = 16'd308;
	#10 start = 1'b1; input_poly1 = 16'd53; input_poly2 = 16'd309;
	#10 start = 1'b1; input_poly1 = 16'd54; input_poly2 = 16'd310;
	#10 start = 1'b1; input_poly1 = 16'd55; input_poly2 = 16'd311;
	#10 start = 1'b1; input_poly1 = 16'd56; input_poly2 = 16'd312;
	#10 start = 1'b1; input_poly1 = 16'd57; input_poly2 = 16'd313;
	#10 start = 1'b1; input_poly1 = 16'd58; input_poly2 = 16'd314;
	#10 start = 1'b1; input_poly1 = 16'd59; input_poly2 = 16'd315;
	#10 start = 1'b1; input_poly1 = 16'd60; input_poly2 = 16'd316;
	#10 start = 1'b1; input_poly1 = 16'd61; input_poly2 = 16'd317;
	#10 start = 1'b1; input_poly1 = 16'd62; input_poly2 = 16'd318;
	#10 start = 1'b1; input_poly1 = 16'd63; input_poly2 = 16'd319;
	#10 start = 1'b1; input_poly1 = 16'd64; input_poly2 = 16'd320;
	#10 start = 1'b1; input_poly1 = 16'd65; input_poly2 = 16'd321;
	#10 start = 1'b1; input_poly1 = 16'd66; input_poly2 = 16'd322;
	#10 start = 1'b1; input_poly1 = 16'd67; input_poly2 = 16'd323;
	#10 start = 1'b1; input_poly1 = 16'd68; input_poly2 = 16'd324;
	#10 start = 1'b1; input_poly1 = 16'd69; input_poly2 = 16'd325;
	#10 start = 1'b1; input_poly1 = 16'd70; input_poly2 = 16'd326;
	#10 start = 1'b1; input_poly1 = 16'd71; input_poly2 = 16'd327;
	#10 start = 1'b1; input_poly1 = 16'd72; input_poly2 = 16'd328;
	#10 start = 1'b1; input_poly1 = 16'd73; input_poly2 = 16'd329;
	#10 start = 1'b1; input_poly1 = 16'd74; input_poly2 = 16'd330;
	#10 start = 1'b1; input_poly1 = 16'd75; input_poly2 = 16'd331;
	#10 start = 1'b1; input_poly1 = 16'd76; input_poly2 = 16'd332;
	#10 start = 1'b1; input_poly1 = 16'd77; input_poly2 = 16'd333;
	#10 start = 1'b1; input_poly1 = 16'd78; input_poly2 = 16'd334;
	#10 start = 1'b1; input_poly1 = 16'd79; input_poly2 = 16'd335;
	#10 start = 1'b1; input_poly1 = 16'd80; input_poly2 = 16'd336;
	#10 start = 1'b1; input_poly1 = 16'd81; input_poly2 = 16'd337;
	#10 start = 1'b1; input_poly1 = 16'd82; input_poly2 = 16'd338;
	#10 start = 1'b1; input_poly1 = 16'd83; input_poly2 = 16'd339;
	#10 start = 1'b1; input_poly1 = 16'd84; input_poly2 = 16'd340;
	#10 start = 1'b1; input_poly1 = 16'd85; input_poly2 = 16'd341;
	#10 start = 1'b1; input_poly1 = 16'd86; input_poly2 = 16'd342;
	#10 start = 1'b1; input_poly1 = 16'd87; input_poly2 = 16'd343;
	#10 start = 1'b1; input_poly1 = 16'd88; input_poly2 = 16'd344;
	#10 start = 1'b1; input_poly1 = 16'd89; input_poly2 = 16'd345;
	#10 start = 1'b1; input_poly1 = 16'd90; input_poly2 = 16'd346;
	#10 start = 1'b1; input_poly1 = 16'd91; input_poly2 = 16'd347;
	#10 start = 1'b1; input_poly1 = 16'd92; input_poly2 = 16'd348;
	#10 start = 1'b1; input_poly1 = 16'd93; input_poly2 = 16'd349;
	#10 start = 1'b1; input_poly1 = 16'd94; input_poly2 = 16'd350;
	#10 start = 1'b1; input_poly1 = 16'd95; input_poly2 = 16'd351;
	#10 start = 1'b1; input_poly1 = 16'd96; input_poly2 = 16'd352;
	#10 start = 1'b1; input_poly1 = 16'd97; input_poly2 = 16'd353;
	#10 start = 1'b1; input_poly1 = 16'd98; input_poly2 = 16'd354;
	#10 start = 1'b1; input_poly1 = 16'd99; input_poly2 = 16'd355;
	#10 start = 1'b1; input_poly1 = 16'd100; input_poly2 = 16'd356;
	#10 start = 1'b1; input_poly1 = 16'd101; input_poly2 = 16'd357;
	#10 start = 1'b1; input_poly1 = 16'd102; input_poly2 = 16'd358;
	#10 start = 1'b1; input_poly1 = 16'd103; input_poly2 = 16'd359;
	#10 start = 1'b1; input_poly1 = 16'd104; input_poly2 = 16'd360;
	#10 start = 1'b1; input_poly1 = 16'd105; input_poly2 = 16'd361;
	#10 start = 1'b1; input_poly1 = 16'd106; input_poly2 = 16'd362;
	#10 start = 1'b1; input_poly1 = 16'd107; input_poly2 = 16'd363;
	#10 start = 1'b1; input_poly1 = 16'd108; input_poly2 = 16'd364;
	#10 start = 1'b1; input_poly1 = 16'd109; input_poly2 = 16'd365;
	#10 start = 1'b1; input_poly1 = 16'd110; input_poly2 = 16'd366;
	#10 start = 1'b1; input_poly1 = 16'd111; input_poly2 = 16'd367;
	#10 start = 1'b1; input_poly1 = 16'd112; input_poly2 = 16'd368;
	#10 start = 1'b1; input_poly1 = 16'd113; input_poly2 = 16'd369;
	#10 start = 1'b1; input_poly1 = 16'd114; input_poly2 = 16'd370;
	#10 start = 1'b1; input_poly1 = 16'd115; input_poly2 = 16'd371;
	#10 start = 1'b1; input_poly1 = 16'd116; input_poly2 = 16'd372;
	#10 start = 1'b1; input_poly1 = 16'd117; input_poly2 = 16'd373;
	#10 start = 1'b1; input_poly1 = 16'd118; input_poly2 = 16'd374;
	#10 start = 1'b1; input_poly1 = 16'd119; input_poly2 = 16'd375;
	#10 start = 1'b1; input_poly1 = 16'd120; input_poly2 = 16'd376;
	#10 start = 1'b1; input_poly1 = 16'd121; input_poly2 = 16'd377;
	#10 start = 1'b1; input_poly1 = 16'd122; input_poly2 = 16'd378;
	#10 start = 1'b1; input_poly1 = 16'd123; input_poly2 = 16'd379;
	#10 start = 1'b1; input_poly1 = 16'd124; input_poly2 = 16'd380;
	#10 start = 1'b1; input_poly1 = 16'd125; input_poly2 = 16'd381;
	#10 start = 1'b1; input_poly1 = 16'd126; input_poly2 = 16'd382;
	#10 start = 1'b1; input_poly1 = 16'd127; input_poly2 = 16'd383;
	#10 start = 1'b1; input_poly1 = 16'd128; input_poly2 = 16'd384;
	#10 start = 1'b1; input_poly1 = 16'd129; input_poly2 = 16'd385;
	#10 start = 1'b1; input_poly1 = 16'd130; input_poly2 = 16'd386;
	#10 start = 1'b1; input_poly1 = 16'd131; input_poly2 = 16'd387;
	#10 start = 1'b1; input_poly1 = 16'd132; input_poly2 = 16'd388;
	#10 start = 1'b1; input_poly1 = 16'd133; input_poly2 = 16'd389;
	#10 start = 1'b1; input_poly1 = 16'd134; input_poly2 = 16'd390;
	#10 start = 1'b1; input_poly1 = 16'd135; input_poly2 = 16'd391;
	#10 start = 1'b1; input_poly1 = 16'd136; input_poly2 = 16'd392;
	#10 start = 1'b1; input_poly1 = 16'd137; input_poly2 = 16'd393;
	#10 start = 1'b1; input_poly1 = 16'd138; input_poly2 = 16'd394;
	#10 start = 1'b1; input_poly1 = 16'd139; input_poly2 = 16'd395;
	#10 start = 1'b1; input_poly1 = 16'd140; input_poly2 = 16'd396;
	#10 start = 1'b1; input_poly1 = 16'd141; input_poly2 = 16'd397;
	#10 start = 1'b1; input_poly1 = 16'd142; input_poly2 = 16'd398;
	#10 start = 1'b1; input_poly1 = 16'd143; input_poly2 = 16'd399;
	#10 start = 1'b1; input_poly1 = 16'd144; input_poly2 = 16'd400;
	#10 start = 1'b1; input_poly1 = 16'd145; input_poly2 = 16'd401;
	#10 start = 1'b1; input_poly1 = 16'd146; input_poly2 = 16'd402;
	#10 start = 1'b1; input_poly1 = 16'd147; input_poly2 = 16'd403;
	#10 start = 1'b1; input_poly1 = 16'd148; input_poly2 = 16'd404;
	#10 start = 1'b1; input_poly1 = 16'd149; input_poly2 = 16'd405;
	#10 start = 1'b1; input_poly1 = 16'd150; input_poly2 = 16'd406;
	#10 start = 1'b1; input_poly1 = 16'd151; input_poly2 = 16'd407;
	#10 start = 1'b1; input_poly1 = 16'd152; input_poly2 = 16'd408;
	#10 start = 1'b1; input_poly1 = 16'd153; input_poly2 = 16'd409;
	#10 start = 1'b1; input_poly1 = 16'd154; input_poly2 = 16'd410;
	#10 start = 1'b1; input_poly1 = 16'd155; input_poly2 = 16'd411;
	#10 start = 1'b1; input_poly1 = 16'd156; input_poly2 = 16'd412;
	#10 start = 1'b1; input_poly1 = 16'd157; input_poly2 = 16'd413;
	#10 start = 1'b1; input_poly1 = 16'd158; input_poly2 = 16'd414;
	#10 start = 1'b1; input_poly1 = 16'd159; input_poly2 = 16'd415;
	#10 start = 1'b1; input_poly1 = 16'd160; input_poly2 = 16'd416;
	#10 start = 1'b1; input_poly1 = 16'd161; input_poly2 = 16'd417;
	#10 start = 1'b1; input_poly1 = 16'd162; input_poly2 = 16'd418;
	#10 start = 1'b1; input_poly1 = 16'd163; input_poly2 = 16'd419;
	#10 start = 1'b1; input_poly1 = 16'd164; input_poly2 = 16'd420;
	#10 start = 1'b1; input_poly1 = 16'd165; input_poly2 = 16'd421;
	#10 start = 1'b1; input_poly1 = 16'd166; input_poly2 = 16'd422;
	#10 start = 1'b1; input_poly1 = 16'd167; input_poly2 = 16'd423;
	#10 start = 1'b1; input_poly1 = 16'd168; input_poly2 = 16'd424;
	#10 start = 1'b1; input_poly1 = 16'd169; input_poly2 = 16'd425;
	#10 start = 1'b1; input_poly1 = 16'd170; input_poly2 = 16'd426;
	#10 start = 1'b1; input_poly1 = 16'd171; input_poly2 = 16'd427;
	#10 start = 1'b1; input_poly1 = 16'd172; input_poly2 = 16'd428;
	#10 start = 1'b1; input_poly1 = 16'd173; input_poly2 = 16'd429;
	#10 start = 1'b1; input_poly1 = 16'd174; input_poly2 = 16'd430;
	#10 start = 1'b1; input_poly1 = 16'd175; input_poly2 = 16'd431;
	#10 start = 1'b1; input_poly1 = 16'd176; input_poly2 = 16'd432;
	#10 start = 1'b1; input_poly1 = 16'd177; input_poly2 = 16'd433;
	#10 start = 1'b1; input_poly1 = 16'd178; input_poly2 = 16'd434;
	#10 start = 1'b1; input_poly1 = 16'd179; input_poly2 = 16'd435;
	#10 start = 1'b1; input_poly1 = 16'd180; input_poly2 = 16'd436;
	#10 start = 1'b1; input_poly1 = 16'd181; input_poly2 = 16'd437;
	#10 start = 1'b1; input_poly1 = 16'd182; input_poly2 = 16'd438;
	#10 start = 1'b1; input_poly1 = 16'd183; input_poly2 = 16'd439;
	#10 start = 1'b1; input_poly1 = 16'd184; input_poly2 = 16'd440;
	#10 start = 1'b1; input_poly1 = 16'd185; input_poly2 = 16'd441;
	#10 start = 1'b1; input_poly1 = 16'd186; input_poly2 = 16'd442;
	#10 start = 1'b1; input_poly1 = 16'd187; input_poly2 = 16'd443;
	#10 start = 1'b1; input_poly1 = 16'd188; input_poly2 = 16'd444;
	#10 start = 1'b1; input_poly1 = 16'd189; input_poly2 = 16'd445;
	#10 start = 1'b1; input_poly1 = 16'd190; input_poly2 = 16'd446;
	#10 start = 1'b1; input_poly1 = 16'd191; input_poly2 = 16'd447;
	#10 start = 1'b1; input_poly1 = 16'd192; input_poly2 = 16'd448;
	#10 start = 1'b1; input_poly1 = 16'd193; input_poly2 = 16'd449;
	#10 start = 1'b1; input_poly1 = 16'd194; input_poly2 = 16'd450;
	#10 start = 1'b1; input_poly1 = 16'd195; input_poly2 = 16'd451;
	#10 start = 1'b1; input_poly1 = 16'd196; input_poly2 = 16'd452;
	#10 start = 1'b1; input_poly1 = 16'd197; input_poly2 = 16'd453;
	#10 start = 1'b1; input_poly1 = 16'd198; input_poly2 = 16'd454;
	#10 start = 1'b1; input_poly1 = 16'd199; input_poly2 = 16'd455;
	#10 start = 1'b1; input_poly1 = 16'd200; input_poly2 = 16'd456;
	#10 start = 1'b1; input_poly1 = 16'd201; input_poly2 = 16'd457;
	#10 start = 1'b1; input_poly1 = 16'd202; input_poly2 = 16'd458;
	#10 start = 1'b1; input_poly1 = 16'd203; input_poly2 = 16'd459;
	#10 start = 1'b1; input_poly1 = 16'd204; input_poly2 = 16'd460;
	#10 start = 1'b1; input_poly1 = 16'd205; input_poly2 = 16'd461;
	#10 start = 1'b1; input_poly1 = 16'd206; input_poly2 = 16'd462;
	#10 start = 1'b1; input_poly1 = 16'd207; input_poly2 = 16'd463;
	#10 start = 1'b1; input_poly1 = 16'd208; input_poly2 = 16'd464;
	#10 start = 1'b1; input_poly1 = 16'd209; input_poly2 = 16'd465;
	#10 start = 1'b1; input_poly1 = 16'd210; input_poly2 = 16'd466;
	#10 start = 1'b1; input_poly1 = 16'd211; input_poly2 = 16'd467;
	#10 start = 1'b1; input_poly1 = 16'd212; input_poly2 = 16'd468;
	#10 start = 1'b1; input_poly1 = 16'd213; input_poly2 = 16'd469;
	#10 start = 1'b1; input_poly1 = 16'd214; input_poly2 = 16'd470;
	#10 start = 1'b1; input_poly1 = 16'd215; input_poly2 = 16'd471;
	#10 start = 1'b1; input_poly1 = 16'd216; input_poly2 = 16'd472;
	#10 start = 1'b1; input_poly1 = 16'd217; input_poly2 = 16'd473;
	#10 start = 1'b1; input_poly1 = 16'd218; input_poly2 = 16'd474;
	#10 start = 1'b1; input_poly1 = 16'd219; input_poly2 = 16'd475;
	#10 start = 1'b1; input_poly1 = 16'd220; input_poly2 = 16'd476;
	#10 start = 1'b1; input_poly1 = 16'd221; input_poly2 = 16'd477;
	#10 start = 1'b1; input_poly1 = 16'd222; input_poly2 = 16'd478;
	#10 start = 1'b1; input_poly1 = 16'd223; input_poly2 = 16'd479;
	#10 start = 1'b1; input_poly1 = 16'd224; input_poly2 = 16'd480;
	#10 start = 1'b1; input_poly1 = 16'd225; input_poly2 = 16'd481;
	#10 start = 1'b1; input_poly1 = 16'd226; input_poly2 = 16'd482;
	#10 start = 1'b1; input_poly1 = 16'd227; input_poly2 = 16'd483;
	#10 start = 1'b1; input_poly1 = 16'd228; input_poly2 = 16'd484;
	#10 start = 1'b1; input_poly1 = 16'd229; input_poly2 = 16'd485;
	#10 start = 1'b1; input_poly1 = 16'd230; input_poly2 = 16'd486;
	#10 start = 1'b1; input_poly1 = 16'd231; input_poly2 = 16'd487;
	#10 start = 1'b1; input_poly1 = 16'd232; input_poly2 = 16'd488;
	#10 start = 1'b1; input_poly1 = 16'd233; input_poly2 = 16'd489;
	#10 start = 1'b1; input_poly1 = 16'd234; input_poly2 = 16'd490;
	#10 start = 1'b1; input_poly1 = 16'd235; input_poly2 = 16'd491;
	#10 start = 1'b1; input_poly1 = 16'd236; input_poly2 = 16'd492;
	#10 start = 1'b1; input_poly1 = 16'd237; input_poly2 = 16'd493;
	#10 start = 1'b1; input_poly1 = 16'd238; input_poly2 = 16'd494;
	#10 start = 1'b1; input_poly1 = 16'd239; input_poly2 = 16'd495;
	#10 start = 1'b1; input_poly1 = 16'd240; input_poly2 = 16'd496;
	#10 start = 1'b1; input_poly1 = 16'd241; input_poly2 = 16'd497;
	#10 start = 1'b1; input_poly1 = 16'd242; input_poly2 = 16'd498;
	#10 start = 1'b1; input_poly1 = 16'd243; input_poly2 = 16'd499;
	#10 start = 1'b1; input_poly1 = 16'd244; input_poly2 = 16'd500;
	#10 start = 1'b1; input_poly1 = 16'd245; input_poly2 = 16'd501;
	#10 start = 1'b1; input_poly1 = 16'd246; input_poly2 = 16'd502;
	#10 start = 1'b1; input_poly1 = 16'd247; input_poly2 = 16'd503;
	#10 start = 1'b1; input_poly1 = 16'd248; input_poly2 = 16'd504;
	#10 start = 1'b1; input_poly1 = 16'd249; input_poly2 = 16'd505;
	#10 start = 1'b1; input_poly1 = 16'd250; input_poly2 = 16'd506;
	#10 start = 1'b1; input_poly1 = 16'd251; input_poly2 = 16'd507;
	#10 start = 1'b1; input_poly1 = 16'd252; input_poly2 = 16'd508;
	#10 start = 1'b1; input_poly1 = 16'd253; input_poly2 = 16'd509;
	#10 start = 1'b1; input_poly1 = 16'd254; input_poly2 = 16'd510;
	#10 start = 1'b1; input_poly1 = 16'd255; input_poly2 = 16'd511;
	#10 start = 1'b1; input_poly1 = 16'd256; input_poly2 = 16'd512;
	#50 start = 1'b0;
	#4000;
	
	#0 start = 1'b0; input_poly1 = 16'd257; input_poly2 = 16'd1;
	#10 start = 1'b1; input_poly1 = 16'd7651; input_poly2 = 16'd1657;
	#10 start = 1'b1; input_poly1 = 16'd3681; input_poly2 = 16'd1026;
	#10 start = 1'b1; input_poly1 = 16'd2503; input_poly2 = 16'd6562;
	#10 start = 1'b1; input_poly1 = 16'd5888; input_poly2 = 16'd4018;
	#10 start = 1'b1; input_poly1 = 16'd505; input_poly2 = 16'd1537;
	#10 start = 1'b1; input_poly1 = 16'd7420; input_poly2 = 16'd6842;
	#10 start = 1'b1; input_poly1 = 16'd3565; input_poly2 = 16'd1289;
	#10 start = 1'b1; input_poly1 = 16'd6133; input_poly2 = 16'd6536;
	#10 start = 1'b1; input_poly1 = 16'd7660; input_poly2 = 16'd1474;
	#10 start = 1'b1; input_poly1 = 16'd7485; input_poly2 = 16'd6399;
	#10 start = 1'b1; input_poly1 = 16'd1027; input_poly2 = 16'd623;
	#10 start = 1'b1; input_poly1 = 16'd4682; input_poly2 = 16'd6885;
	#10 start = 1'b1; input_poly1 = 16'd1870; input_poly2 = 16'd7127;
	#10 start = 1'b1; input_poly1 = 16'd4366; input_poly2 = 16'd703;
	#10 start = 1'b1; input_poly1 = 16'd1706; input_poly2 = 16'd1981;
	#10 start = 1'b1; input_poly1 = 16'd6463; input_poly2 = 16'd406;
	#10 start = 1'b1; input_poly1 = 16'd2247; input_poly2 = 16'd1172;
	#10 start = 1'b1; input_poly1 = 16'd5457; input_poly2 = 16'd5683;
	#10 start = 1'b1; input_poly1 = 16'd5126; input_poly2 = 16'd5434;
	#10 start = 1'b1; input_poly1 = 16'd1215; input_poly2 = 16'd7082;
	#10 start = 1'b1; input_poly1 = 16'd6834; input_poly2 = 16'd780;
	#10 start = 1'b1; input_poly1 = 16'd2784; input_poly2 = 16'd2473;
	#10 start = 1'b1; input_poly1 = 16'd7472; input_poly2 = 16'd6043;
	#10 start = 1'b1; input_poly1 = 16'd850; input_poly2 = 16'd6550;
	#10 start = 1'b1; input_poly1 = 16'd7608; input_poly2 = 16'd3124;
	#10 start = 1'b1; input_poly1 = 16'd3196; input_poly2 = 16'd6424;
	#10 start = 1'b1; input_poly1 = 16'd519; input_poly2 = 16'd5309;
	#10 start = 1'b1; input_poly1 = 16'd2032; input_poly2 = 16'd5345;
	#10 start = 1'b1; input_poly1 = 16'd3420; input_poly2 = 16'd4279;
	#10 start = 1'b1; input_poly1 = 16'd4209; input_poly2 = 16'd7218;
	#10 start = 1'b1; input_poly1 = 16'd6082; input_poly2 = 16'd5196;
	#10 start = 1'b1; input_poly1 = 16'd4295; input_poly2 = 16'd5583;
	#10 start = 1'b1; input_poly1 = 16'd1383; input_poly2 = 16'd1174;
	#10 start = 1'b1; input_poly1 = 16'd1761; input_poly2 = 16'd7321;
	#10 start = 1'b1; input_poly1 = 16'd5951; input_poly2 = 16'd5444;
	#10 start = 1'b1; input_poly1 = 16'd5660; input_poly2 = 16'd5844;
	#10 start = 1'b1; input_poly1 = 16'd457; input_poly2 = 16'd6970;
	#10 start = 1'b1; input_poly1 = 16'd6357; input_poly2 = 16'd5690;
	#10 start = 1'b1; input_poly1 = 16'd7374; input_poly2 = 16'd6530;
	#10 start = 1'b1; input_poly1 = 16'd4244; input_poly2 = 16'd5996;
	#10 start = 1'b1; input_poly1 = 16'd1950; input_poly2 = 16'd7587;
	#10 start = 1'b1; input_poly1 = 16'd2333; input_poly2 = 16'd4946;
	#10 start = 1'b1; input_poly1 = 16'd1625; input_poly2 = 16'd753;
	#10 start = 1'b1; input_poly1 = 16'd4914; input_poly2 = 16'd743;
	#10 start = 1'b1; input_poly1 = 16'd2334; input_poly2 = 16'd2476;
	#10 start = 1'b1; input_poly1 = 16'd4831; input_poly2 = 16'd5871;
	#10 start = 1'b1; input_poly1 = 16'd4406; input_poly2 = 16'd4005;
	#10 start = 1'b1; input_poly1 = 16'd2700; input_poly2 = 16'd7564;
	#10 start = 1'b1; input_poly1 = 16'd7441; input_poly2 = 16'd5696;
	#10 start = 1'b1; input_poly1 = 16'd1132; input_poly2 = 16'd4700;
	#10 start = 1'b1; input_poly1 = 16'd3416; input_poly2 = 16'd1120;
	#10 start = 1'b1; input_poly1 = 16'd3719; input_poly2 = 16'd4737;
	#10 start = 1'b1; input_poly1 = 16'd3751; input_poly2 = 16'd5429;
	#10 start = 1'b1; input_poly1 = 16'd6140; input_poly2 = 16'd6978;
	#10 start = 1'b1; input_poly1 = 16'd4201; input_poly2 = 16'd3846;
	#10 start = 1'b1; input_poly1 = 16'd4935; input_poly2 = 16'd1411;
	#10 start = 1'b1; input_poly1 = 16'd6717; input_poly2 = 16'd3875;
	#10 start = 1'b1; input_poly1 = 16'd882; input_poly2 = 16'd5829;
	#10 start = 1'b1; input_poly1 = 16'd3018; input_poly2 = 16'd4729;
	#10 start = 1'b1; input_poly1 = 16'd3051; input_poly2 = 16'd6470;
	#10 start = 1'b1; input_poly1 = 16'd6976; input_poly2 = 16'd5659;
	#10 start = 1'b1; input_poly1 = 16'd638; input_poly2 = 16'd2574;
	#10 start = 1'b1; input_poly1 = 16'd7058; input_poly2 = 16'd4742;
	#10 start = 1'b1; input_poly1 = 16'd1298; input_poly2 = 16'd4952;
	#10 start = 1'b1; input_poly1 = 16'd2367; input_poly2 = 16'd6462;
	#10 start = 1'b1; input_poly1 = 16'd6131; input_poly2 = 16'd3183;
	#10 start = 1'b1; input_poly1 = 16'd2327; input_poly2 = 16'd667;
	#10 start = 1'b1; input_poly1 = 16'd507; input_poly2 = 16'd4363;
	#10 start = 1'b1; input_poly1 = 16'd5265; input_poly2 = 16'd1668;
	#10 start = 1'b1; input_poly1 = 16'd1854; input_poly2 = 16'd2469;
	#10 start = 1'b1; input_poly1 = 16'd5522; input_poly2 = 16'd4044;
	#10 start = 1'b1; input_poly1 = 16'd3025; input_poly2 = 16'd2358;
	#10 start = 1'b1; input_poly1 = 16'd7123; input_poly2 = 16'd418;
	#10 start = 1'b1; input_poly1 = 16'd2530; input_poly2 = 16'd6834;
	#10 start = 1'b1; input_poly1 = 16'd1668; input_poly2 = 16'd2754;
	#10 start = 1'b1; input_poly1 = 16'd838; input_poly2 = 16'd5218;
	#10 start = 1'b1; input_poly1 = 16'd2169; input_poly2 = 16'd5979;
	#10 start = 1'b1; input_poly1 = 16'd4196; input_poly2 = 16'd1061;
	#10 start = 1'b1; input_poly1 = 16'd3015; input_poly2 = 16'd3487;
	#10 start = 1'b1; input_poly1 = 16'd7369; input_poly2 = 16'd5669;
	#10 start = 1'b1; input_poly1 = 16'd7219; input_poly2 = 16'd3984;
	#10 start = 1'b1; input_poly1 = 16'd6934; input_poly2 = 16'd1299;
	#10 start = 1'b1; input_poly1 = 16'd4589; input_poly2 = 16'd7218;
	#10 start = 1'b1; input_poly1 = 16'd2842; input_poly2 = 16'd3783;
	#10 start = 1'b1; input_poly1 = 16'd6537; input_poly2 = 16'd4171;
	#10 start = 1'b1; input_poly1 = 16'd3890; input_poly2 = 16'd5010;
	#10 start = 1'b1; input_poly1 = 16'd282; input_poly2 = 16'd4287;
	#10 start = 1'b1; input_poly1 = 16'd3080; input_poly2 = 16'd6334;
	#10 start = 1'b1; input_poly1 = 16'd7494; input_poly2 = 16'd5894;
	#10 start = 1'b1; input_poly1 = 16'd4180; input_poly2 = 16'd7398;
	#10 start = 1'b1; input_poly1 = 16'd3533; input_poly2 = 16'd4564;
	#10 start = 1'b1; input_poly1 = 16'd6969; input_poly2 = 16'd1623;
	#10 start = 1'b1; input_poly1 = 16'd3741; input_poly2 = 16'd3192;
	#10 start = 1'b1; input_poly1 = 16'd2439; input_poly2 = 16'd7626;
	#10 start = 1'b1; input_poly1 = 16'd2720; input_poly2 = 16'd4057;
	#10 start = 1'b1; input_poly1 = 16'd1961; input_poly2 = 16'd2189;
	#10 start = 1'b1; input_poly1 = 16'd2260; input_poly2 = 16'd5378;
	#10 start = 1'b1; input_poly1 = 16'd4978; input_poly2 = 16'd2086;
	#10 start = 1'b1; input_poly1 = 16'd1562; input_poly2 = 16'd1908;
	#10 start = 1'b1; input_poly1 = 16'd6879; input_poly2 = 16'd4140;
	#10 start = 1'b1; input_poly1 = 16'd951; input_poly2 = 16'd3022;
	#10 start = 1'b1; input_poly1 = 16'd6467; input_poly2 = 16'd3096;
	#10 start = 1'b1; input_poly1 = 16'd5821; input_poly2 = 16'd4497;
	#10 start = 1'b1; input_poly1 = 16'd2484; input_poly2 = 16'd3822;
	#10 start = 1'b1; input_poly1 = 16'd1363; input_poly2 = 16'd4549;
	#10 start = 1'b1; input_poly1 = 16'd1234; input_poly2 = 16'd2713;
	#10 start = 1'b1; input_poly1 = 16'd5950; input_poly2 = 16'd4591;
	#10 start = 1'b1; input_poly1 = 16'd4090; input_poly2 = 16'd7621;
	#10 start = 1'b1; input_poly1 = 16'd3097; input_poly2 = 16'd6860;
	#10 start = 1'b1; input_poly1 = 16'd5725; input_poly2 = 16'd1126;
	#10 start = 1'b1; input_poly1 = 16'd2914; input_poly2 = 16'd3853;
	#10 start = 1'b1; input_poly1 = 16'd6284; input_poly2 = 16'd6946;
	#10 start = 1'b1; input_poly1 = 16'd1720; input_poly2 = 16'd2369;
	#10 start = 1'b1; input_poly1 = 16'd6933; input_poly2 = 16'd2804;
	#10 start = 1'b1; input_poly1 = 16'd5318; input_poly2 = 16'd6984;
	#10 start = 1'b1; input_poly1 = 16'd1040; input_poly2 = 16'd2873;
	#10 start = 1'b1; input_poly1 = 16'd2089; input_poly2 = 16'd7399;
	#10 start = 1'b1; input_poly1 = 16'd584; input_poly2 = 16'd3430;
	#10 start = 1'b1; input_poly1 = 16'd6908; input_poly2 = 16'd1451;
	#10 start = 1'b1; input_poly1 = 16'd1916; input_poly2 = 16'd3300;
	#10 start = 1'b1; input_poly1 = 16'd618; input_poly2 = 16'd2376;
	#10 start = 1'b1; input_poly1 = 16'd3171; input_poly2 = 16'd3139;
	#10 start = 1'b1; input_poly1 = 16'd1712; input_poly2 = 16'd341;
	#10 start = 1'b1; input_poly1 = 16'd5939; input_poly2 = 16'd4795;
	#10 start = 1'b1; input_poly1 = 16'd2350; input_poly2 = 16'd7304;
	#10 start = 1'b1; input_poly1 = 16'd7219; input_poly2 = 16'd786;
	#10 start = 1'b1; input_poly1 = 16'd6689; input_poly2 = 16'd4036;
	#10 start = 1'b1; input_poly1 = 16'd7475; input_poly2 = 16'd6140;
	#10 start = 1'b1; input_poly1 = 16'd1527; input_poly2 = 16'd6543;
	#10 start = 1'b1; input_poly1 = 16'd340; input_poly2 = 16'd299;
	#10 start = 1'b1; input_poly1 = 16'd451; input_poly2 = 16'd2345;
	#10 start = 1'b1; input_poly1 = 16'd1095; input_poly2 = 16'd7534;
	#10 start = 1'b1; input_poly1 = 16'd402; input_poly2 = 16'd7183;
	#10 start = 1'b1; input_poly1 = 16'd2620; input_poly2 = 16'd7240;
	#10 start = 1'b1; input_poly1 = 16'd3438; input_poly2 = 16'd6399;
	#10 start = 1'b1; input_poly1 = 16'd7026; input_poly2 = 16'd590;
	#10 start = 1'b1; input_poly1 = 16'd6973; input_poly2 = 16'd7083;
	#10 start = 1'b1; input_poly1 = 16'd588; input_poly2 = 16'd1004;
	#10 start = 1'b1; input_poly1 = 16'd5242; input_poly2 = 16'd5532;
	#10 start = 1'b1; input_poly1 = 16'd1726; input_poly2 = 16'd4156;
	#10 start = 1'b1; input_poly1 = 16'd7422; input_poly2 = 16'd332;
	#10 start = 1'b1; input_poly1 = 16'd5500; input_poly2 = 16'd1423;
	#10 start = 1'b1; input_poly1 = 16'd4884; input_poly2 = 16'd400;
	#10 start = 1'b1; input_poly1 = 16'd6434; input_poly2 = 16'd3992;
	#10 start = 1'b1; input_poly1 = 16'd1770; input_poly2 = 16'd1430;
	#10 start = 1'b1; input_poly1 = 16'd6527; input_poly2 = 16'd2606;
	#10 start = 1'b1; input_poly1 = 16'd4813; input_poly2 = 16'd1984;
	#10 start = 1'b1; input_poly1 = 16'd3650; input_poly2 = 16'd5957;
	#10 start = 1'b1; input_poly1 = 16'd7295; input_poly2 = 16'd3559;
	#10 start = 1'b1; input_poly1 = 16'd1521; input_poly2 = 16'd3825;
	#10 start = 1'b1; input_poly1 = 16'd6121; input_poly2 = 16'd669;
	#10 start = 1'b1; input_poly1 = 16'd1360; input_poly2 = 16'd2377;
	#10 start = 1'b1; input_poly1 = 16'd6800; input_poly2 = 16'd5614;
	#10 start = 1'b1; input_poly1 = 16'd4320; input_poly2 = 16'd1870;
	#10 start = 1'b1; input_poly1 = 16'd1096; input_poly2 = 16'd5329;
	#10 start = 1'b1; input_poly1 = 16'd3417; input_poly2 = 16'd3873;
	#10 start = 1'b1; input_poly1 = 16'd1103; input_poly2 = 16'd3148;
	#10 start = 1'b1; input_poly1 = 16'd2484; input_poly2 = 16'd5356;
	#10 start = 1'b1; input_poly1 = 16'd1519; input_poly2 = 16'd5800;
	#10 start = 1'b1; input_poly1 = 16'd3426; input_poly2 = 16'd1348;
	#10 start = 1'b1; input_poly1 = 16'd2217; input_poly2 = 16'd664;
	#10 start = 1'b1; input_poly1 = 16'd4808; input_poly2 = 16'd1312;
	#10 start = 1'b1; input_poly1 = 16'd3308; input_poly2 = 16'd7106;
	#10 start = 1'b1; input_poly1 = 16'd5222; input_poly2 = 16'd5920;
	#10 start = 1'b1; input_poly1 = 16'd5320; input_poly2 = 16'd2706;
	#10 start = 1'b1; input_poly1 = 16'd828; input_poly2 = 16'd2759;
	#10 start = 1'b1; input_poly1 = 16'd2041; input_poly2 = 16'd7284;
	#10 start = 1'b1; input_poly1 = 16'd6343; input_poly2 = 16'd3183;
	#10 start = 1'b1; input_poly1 = 16'd7654; input_poly2 = 16'd1418;
	#10 start = 1'b1; input_poly1 = 16'd3354; input_poly2 = 16'd6051;
	#10 start = 1'b1; input_poly1 = 16'd1949; input_poly2 = 16'd5640;
	#10 start = 1'b1; input_poly1 = 16'd7076; input_poly2 = 16'd620;
	#10 start = 1'b1; input_poly1 = 16'd5936; input_poly2 = 16'd3086;
	#10 start = 1'b1; input_poly1 = 16'd1558; input_poly2 = 16'd360;
	#10 start = 1'b1; input_poly1 = 16'd6888; input_poly2 = 16'd3564;
	#10 start = 1'b1; input_poly1 = 16'd7251; input_poly2 = 16'd1008;
	#10 start = 1'b1; input_poly1 = 16'd6039; input_poly2 = 16'd1826;
	#10 start = 1'b1; input_poly1 = 16'd4111; input_poly2 = 16'd2616;
	#10 start = 1'b1; input_poly1 = 16'd2287; input_poly2 = 16'd7653;
	#10 start = 1'b1; input_poly1 = 16'd2433; input_poly2 = 16'd7236;
	#10 start = 1'b1; input_poly1 = 16'd4283; input_poly2 = 16'd6296;
	#10 start = 1'b1; input_poly1 = 16'd3633; input_poly2 = 16'd2688;
	#10 start = 1'b1; input_poly1 = 16'd701; input_poly2 = 16'd5966;
	#10 start = 1'b1; input_poly1 = 16'd5149; input_poly2 = 16'd7332;
	#10 start = 1'b1; input_poly1 = 16'd4576; input_poly2 = 16'd6697;
	#10 start = 1'b1; input_poly1 = 16'd1522; input_poly2 = 16'd2114;
	#10 start = 1'b1; input_poly1 = 16'd5516; input_poly2 = 16'd4650;
	#10 start = 1'b1; input_poly1 = 16'd2249; input_poly2 = 16'd1581;
	#10 start = 1'b1; input_poly1 = 16'd2679; input_poly2 = 16'd3329;
	#10 start = 1'b1; input_poly1 = 16'd7061; input_poly2 = 16'd3469;
	#10 start = 1'b1; input_poly1 = 16'd1634; input_poly2 = 16'd711;
	#10 start = 1'b1; input_poly1 = 16'd3077; input_poly2 = 16'd4426;
	#10 start = 1'b1; input_poly1 = 16'd4935; input_poly2 = 16'd433;
	#10 start = 1'b1; input_poly1 = 16'd283; input_poly2 = 16'd995;
	#10 start = 1'b1; input_poly1 = 16'd3378; input_poly2 = 16'd6496;
	#10 start = 1'b1; input_poly1 = 16'd6411; input_poly2 = 16'd4364;
	#10 start = 1'b1; input_poly1 = 16'd2228; input_poly2 = 16'd5363;
	#10 start = 1'b1; input_poly1 = 16'd2328; input_poly2 = 16'd7307;
	#10 start = 1'b1; input_poly1 = 16'd7303; input_poly2 = 16'd1280;
	#10 start = 1'b1; input_poly1 = 16'd5866; input_poly2 = 16'd3435;
	#10 start = 1'b1; input_poly1 = 16'd7322; input_poly2 = 16'd3185;
	#10 start = 1'b1; input_poly1 = 16'd6698; input_poly2 = 16'd2718;
	#10 start = 1'b1; input_poly1 = 16'd6596; input_poly2 = 16'd4593;
	#10 start = 1'b1; input_poly1 = 16'd3159; input_poly2 = 16'd6807;
	#10 start = 1'b1; input_poly1 = 16'd1270; input_poly2 = 16'd6535;
	#10 start = 1'b1; input_poly1 = 16'd2607; input_poly2 = 16'd4074;
	#10 start = 1'b1; input_poly1 = 16'd1616; input_poly2 = 16'd3997;
	#10 start = 1'b1; input_poly1 = 16'd2653; input_poly2 = 16'd3276;
	#10 start = 1'b1; input_poly1 = 16'd4797; input_poly2 = 16'd4130;
	#10 start = 1'b1; input_poly1 = 16'd3651; input_poly2 = 16'd6685;
	#10 start = 1'b1; input_poly1 = 16'd4865; input_poly2 = 16'd1307;
	#10 start = 1'b1; input_poly1 = 16'd6224; input_poly2 = 16'd4228;
	#10 start = 1'b1; input_poly1 = 16'd6250; input_poly2 = 16'd1031;
	#10 start = 1'b1; input_poly1 = 16'd4301; input_poly2 = 16'd4512;
	#10 start = 1'b1; input_poly1 = 16'd4461; input_poly2 = 16'd1788;
	#10 start = 1'b1; input_poly1 = 16'd2651; input_poly2 = 16'd3405;
	#10 start = 1'b1; input_poly1 = 16'd5926; input_poly2 = 16'd4644;
	#10 start = 1'b1; input_poly1 = 16'd2643; input_poly2 = 16'd3097;
	#10 start = 1'b1; input_poly1 = 16'd5075; input_poly2 = 16'd3161;
	#10 start = 1'b1; input_poly1 = 16'd2741; input_poly2 = 16'd7513;
	#10 start = 1'b1; input_poly1 = 16'd2587; input_poly2 = 16'd6375;
	#10 start = 1'b1; input_poly1 = 16'd2978; input_poly2 = 16'd4309;
	#10 start = 1'b1; input_poly1 = 16'd5075; input_poly2 = 16'd327;
	#10 start = 1'b1; input_poly1 = 16'd3500; input_poly2 = 16'd2572;
	#10 start = 1'b1; input_poly1 = 16'd3460; input_poly2 = 16'd4044;
	#10 start = 1'b1; input_poly1 = 16'd1128; input_poly2 = 16'd1054;
	#10 start = 1'b1; input_poly1 = 16'd5395; input_poly2 = 16'd4426;
	#10 start = 1'b1; input_poly1 = 16'd5498; input_poly2 = 16'd2476;
	#10 start = 1'b1; input_poly1 = 16'd754; input_poly2 = 16'd2151;
	#10 start = 1'b1; input_poly1 = 16'd7322; input_poly2 = 16'd4707;
	#10 start = 1'b1; input_poly1 = 16'd1106; input_poly2 = 16'd3738;
	#10 start = 1'b1; input_poly1 = 16'd7528; input_poly2 = 16'd6497;
	#10 start = 1'b1; input_poly1 = 16'd1596; input_poly2 = 16'd2928;
	#10 start = 1'b1; input_poly1 = 16'd6386; input_poly2 = 16'd4583;
	#10 start = 1'b1; input_poly1 = 16'd2873; input_poly2 = 16'd2404;
	#10 start = 1'b1; input_poly1 = 16'd4103; input_poly2 = 16'd7097;
	#10 start = 1'b1; input_poly1 = 16'd1802; input_poly2 = 16'd7608;
	#10 start = 1'b1; input_poly1 = 16'd7654; input_poly2 = 16'd4057;
	#10 start = 1'b1; input_poly1 = 16'd6801; input_poly2 = 16'd3609;
	#10 start = 1'b1; input_poly1 = 16'd3981; input_poly2 = 16'd1759;
	#10 start = 1'b1; input_poly1 = 16'd5404; input_poly2 = 16'd1646;
	#10 start = 1'b1; input_poly1 = 16'd3881; input_poly2 = 16'd517;
	#10 start = 1'b1; input_poly1 = 16'd5318; input_poly2 = 16'd7416;
	#10 start = 1'b1; input_poly1 = 16'd3049; input_poly2 = 16'd5444;
	#10 start = 1'b1; input_poly1 = 16'd3833; input_poly2 = 16'd979;
	#10 start = 1'b1; input_poly1 = 16'd5194; input_poly2 = 16'd4540;
	#10 start = 1'b1; input_poly1 = 16'd4940; input_poly2 = 16'd7549;
	#10 start = 1'b1; input_poly1 = 16'd1590; input_poly2 = 16'd6913;
	#10 start = 1'b1; input_poly1 = 16'd4234; input_poly2 = 16'd5215;
	#10 start = 1'b1; input_poly1 = 16'd2771; input_poly2 = 16'd1326;
	#10 start = 1'b1; input_poly1 = 16'd6575; input_poly2 = 16'd3488;
	#10 start = 1'b1; input_poly1 = 16'd336; input_poly2 = 16'd2766;
	#10 start = 1'b1; input_poly1 = 16'd3050; input_poly2 = 16'd1401;
	#10 start = 1'b1; input_poly1 = 16'd4519; input_poly2 = 16'd5142;
	#10 start = 1'b1; input_poly1 = 16'd6274; input_poly2 = 16'd7203;
	#10 start = 1'b1; input_poly1 = 16'd4518; input_poly2 = 16'd3505;
	#50 start = 1'b0;
	
	
	#6000 $stop;
	
	end
    
    
endmodule
